module prop ();
   wire prop;
endmodule

