// Author: Aman Goel (amangoel@umich.edu), University of Michigan

module prop ();
   wire prop;
endmodule

